CIRCUIT C:\Documents and Settings\Administrator\My Documents\microwind3\Book mw CMOS\inv.MSK
*
* IC Technology: CMOS 0.12�m - 6 Metal
*
VDD 1 0 DC 1.20
Vin 6 0 PULSE(0.00 1.20 0.23N 0.02N 0.02N 0.23N 0.50N)
*
* List of nodes
* "inv" corresponds to n�3
* "N5" corresponds to n�5
* "in" corresponds to n�6
* "N7" corresponds to n�7
*
* MOS devices
MN1 0 6 3 0 N1  W= 0.24U L= 0.12U
MP1 1 6 3 1 P1  W= 0.72U L= 0.12U
*
C2 1 0  1.340fF
C3 3 0  1.033fF
C5 5 0  0.080fF
C6 6 0  0.314fF
C7 7 0  0.035fF
*
* n-MOS Model 3 :
* low leakage
.MODEL N1 NMOS LEVEL=3 VTO=0.40 UO=600.000 TOX= 2.0E-9
+LD =0.000U THETA=0.500 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=120.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* p-MOS Model 3:
* low leakage
.MODEL P1 PMOS LEVEL=3 VTO=-0.45 UO=200.000 TOX= 2.0E-9
+LD =0.000U THETA=0.300 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=110.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* Transient analysis
*
.TEMP 27.0
.TRAN 0.1N 2.00N
* (Pspice)
.PROBE
.END
